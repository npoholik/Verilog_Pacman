`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/20/2025 03:12:38 PM
// Design Name: 
// Module Name: Pac_Sprite
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//  
//////////////////////////////////////////////////////////////////////////////////

module Map_Access (
    input signed [10:0] x_VGA, y_VGA, 
    output reg [5:0] GRID_TYPE          // Accessing the type of grid on the map
);

//**** DEFINE MAP GRID *** //
// Need to define macros (not all might be used):
localparam BLNK = 0;
localparam BVWE = 1 /* Border vertical wall*/; localparam BVWW = 2; localparam BHWN = 3; localparam BHWS = 4 /* Border horizontal wall*/;
localparam BCNE = 5 /* border corner north to east*/; localparam BCES = 6; localparam BCSW = 7; localparam BCWN = 8;
localparam BTWE = 9 /* border T wall east*/; localparam BTWW = 10; localparam BTWN = 11; localparam BTWS = 12; 
localparam SCNE = 13 /* shallow corner north to east*/; localparam SCES = 14; localparam SCSW = 15; localparam SCWN = 16; 
localparam DCNE = 17 /* deep corner north to east */; localparam DCES = 18; localparam DCSW = 19; localparam DCWN = 20;
localparam IMWW = 21 /* Interior map wall west */; localparam IMWE = 22; localparam IMWN = 23; localparam IMWS = 24; 
localparam MMGG = 25 /*map middle ghost gate */; 

logic [11:0] gridMap [0:27][0:35] = '{
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK}, 
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK},
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK},
    '{BCNE, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BTWW, BTWE, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BHWN, BCES}, 
    '{BVWW, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BVWE}, 
    '{BVWW, BLNK, SCNE, IMWN, IMWN, SCES, BLNK, SCNE, IMWN, IMWN, IMWN, SCES, BLNK, IMWW, IMWE, BLNK, SCNE, IMWN, IMWN, IMWN, SCES, BLNK, SCNE, IMWN, IMWN, SCES, BLNK, BVWE}, 
    '{BVWW, BLNK, IMWW, BLNK, BLNK, IMWE, BLNK, IMWW, BLNK, BLNK, BLNK, IMWE, BLNK, IMWW, IMWE, BLNK, IMWW, BLNK, BLNK, BLNK, IMWE, BLNK, IMWW, BLNK, BLNK, IMWE, BLNK, BVWE}, 
    '{BVWW, BLNK, SCWN, IMWS, IMWS, SCSW, BLNK, SCWN, IMWS, IMWS, IMWS, SCSW, BLNK, SCWN, SCSW, BLNK, SCWN, IMWS, IMWS, IMWS, SCSW, BLNK, SCWN, IMWS, IMWS, SCSW, BLNK, BVWE}, 
    '{BVWW, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BVWE}, 
    '{BVWW, BLNK, SCNE, IMWN, IMWN, SCES, BLNK, SCNE, SCES, BLNK, SCNE, IMWN, IMWN, IMWN, IMWN, IMWN, IMWN, SCES, BLNK, SCNE, SCES, BLNK, SCNE, IMWN, IMWN, SCES, BLNK, BVWE}, 
    '{BVWW, BLNK, SCWN, IMWS, IMWS, SCSW, BLNK, IMWW, IMWE, BLNK, SCWN, IMWS, IMWS, DCES, DCNE, IMWS, IMWS, SCSW, BLNK, IMWW, IMWE, BLNK, SCWN, IMWS, IMWS, SCSW, BLNK, BVWE}, 
    '{BVWW, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BVWE}, 
    '{BCWN, BHWS, BHWS, BHWS, BHWS, SCES, BLNK, IMWW, DCWN, IMWN, IMWN, SCES, BLNK, IMWW, IMWE, BLNK, SCNE, IMWN, IMWN, DCSW, IMWE, BLNK, SCNE, BHWS, BHWS, BHWS, BHWS, BCSW}, 
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BVWW, BLNK, IMWW, DCNE, IMWS, IMWS, SCSW, BLNK, SCWN, SCSW, BLNK, SCWN, IMWS, IMWS, DCES, IMWE, BLNK, BVWE, BLNK, BLNK, BLNK, BLNK, BLNK}, 
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BVWW, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BVWE, BLNK, BLNK, BLNK, BLNK, BLNK}, 
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BVWW, BLNK, IMWW, IMWE, BLNK, SCNE, IMWN, IMWN, MMGG, MMGG, IMWN, IMWN, SCES, BLNK, IMWW, IMWE, BLNK, BVWE, BLNK, BLNK, BLNK, BLNK, BLNK}, 
    '{BHWN, BHWN, BHWN, BHWN, BHWN, SCSW, BLNK, SCWN, SCSW, BLNK, IMWW, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWE, BLNK, SCWN, SCSW, BLNK, SCWN, BHWN, BHWN, BHWN, BHWN, BHWN}, 
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWW, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWE, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK}, 
    '{BHWS, BHWS, BHWS, BHWS, BHWS, SCES, BLNK, SCNE, SCES, BLNK, IMWW, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWE, BLNK, SCNE, SCES, BLNK, SCNE, BHWS, BHWS, BHWS, BHWS, BHWS}, 
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BVWW, BLNK, IMWW, IMWE, BLNK, SCWN, IMWS, IMWS, IMWS, IMWS, IMWS, IMWS, SCSW, BLNK, IMWW, IMWE, BLNK, BVWE, BLNK, BLNK, BLNK, BLNK, BLNK}, 
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BVWW, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BVWE, BLNK, BLNK, BLNK, BLNK, BLNK}, 
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BVWW, BLNK, IMWW, IMWE, BLNK, SCNE, IMWN, IMWN, IMWN, IMWN, IMWN, IMWN, SCES, BLNK, IMWW, IMWE, BLNK, BVWE, BLNK, BLNK, BLNK, BLNK, BLNK}, 
    '{BCNE, BHWN, BHWN, BHWN, BHWN, SCSW, BLNK, SCWN, SCSW, BLNK, SCWN, IMWS, IMWS, DCES, DCNE, IMWS, IMWS, SCSW, BLNK, SCWN, SCSW, BLNK, SCWN, BHWN, BHWN, BHWN, BHWN, BCES}, 
    '{BVWW, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BVWE}, 
    '{BVWW, BLNK, SCNE, IMWN, IMWN, SCES, BLNK, SCNE, IMWN, IMWN, IMWN, SCES, BLNK, IMWW, IMWE, BLNK, SCNE, IMWN, IMWN, IMWN, SCES, BLNK, SCNE, IMWN, IMWN, SCES, BLNK, BVWE}, 
    '{BVWW, BLNK, SCWN, IMWS, DCES, IMWE, BLNK, SCWN, IMWS, IMWS, IMWS, SCSW, BLNK, SCWN, SCSW, BLNK, SCWN, IMWS, IMWS, IMWS, SCSW, BLNK, IMWW, DCNE, IMWS, SCSW, BLNK, BVWE}, 
    '{BVWW, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BVWE}, 
    '{BTWN, IMWN, SCES, BLNK, IMWW, IMWE, BLNK, SCNE, SCES, BLNK, SCNE, IMWN, IMWN, IMWN, IMWN, IMWN, IMWN, SCES, BLNK, SCNE, SCES, BLNK, IMWW, IMWE, BLNK, SCNE, IMWN, BTWN}, 
    '{BTWS, IMWS, SCSW, BLNK, SCWN, SCSW, BLNK, IMWW, IMWE, BLNK, SCWN, IMWS, IMWS, DCES, DCNE, IMWS, IMWS, SCSW, BLNK, IMWW, IMWE, BLNK, SCWN, SCSW, BLNK, SCWN, IMWS, BTWS}, 
    '{BVWW, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, IMWW, IMWE, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BVWE}, 
    '{BVWW, BLNK, SCNE, IMWN, IMWN, IMWN, IMWN, DCSW, DCWN, IMWN, IMWN, SCES, BLNK, IMWW, IMWE, BLNK, SCNE, IMWN, IMWN, DCSW, DCWN, IMWN, IMWN, IMWN, IMWN, SCES, BLNK, BVWE}, 
    '{BVWW, BLNK, SCWN, IMWS, IMWS, IMWS, IMWS, IMWS, IMWS, IMWS, IMWS, SCSW, BLNK, SCWN, SCSW, BLNK, SCWN, IMWS, IMWS, IMWS, IMWS, IMWS, IMWS, IMWS, IMWS, SCSW, BLNK, BVWE}, 
    '{BVWW, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BVWE}, 
    '{BCWN, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BHWS, BCSW}, 
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK},
    '{BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK, BLNK} };

endmodule 
